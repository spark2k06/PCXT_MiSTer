`ifndef KF8255_DEFINITIONS_SVH
`define KF8255_DEFINITIONS_SVH

`define ADDRESS_PORT_A          (2'b00)
`define ADDRESS_PORT_B          (2'b01)
`define ADDRESS_PORT_C          (2'b10)
`define ADDRESS_CONTROL         (2'b11)

`define KF8255_CONTROL_MODE_0   (2'b00)
`define KF8255_CONTROL_MODE_1   (2'b01)
`define KF8255_CONTROL_MODE_2   (2'b1?)

`define PORT_INPUT              (1'b1)
`define PORT_OUTPUT             (1'b0)

`endif
